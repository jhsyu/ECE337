// $Id: $
// File name:   tb_mealy.sv
// Created:     9/29/2020
// Author:      Jiahao Xu
// Lab Section: 337-002
// Version:     1.0  Initial Design Entry
// Description: . 

module tb_mealy ();

endmodule