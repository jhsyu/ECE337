// $Id: $
// File name:   ahb_lite_fir_filter.sv
// Created:     10/27/2020
// Author:      Jiahao Xu
// Lab Section: 337-002
// Version:     1.0  Initial Design Entry
// Description: . 
